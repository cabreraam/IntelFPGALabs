module char_7seg_hex (C, Display);

  input [3:0] C;
  output [6:0] Display;

  assign Display =
    (C == 4'b0000) ? 7'b1000000 : // 0
    (C == 4'b0001) ? 7'b1111001 : // 1
    (C == 4'b0010) ? 7'b0100100 : // 2
    (C == 4'b0011) ? 7'b0110000 : // 3
    (C == 4'b0100) ? 7'b0011001 : // 4
    (C == 4'b0101) ? 7'b0010010 : // 5
    (C == 4'b0110) ? 7'b0000010 : // 6
    (C == 4'b0111) ? 7'b1111000 : // 7
    (C == 4'b1000) ? 7'b0000000 : // 8
    (C == 4'b1001) ? 7'b0011000 : // 9
    (C == 4'b1010) ? 7'b0001000 : // a
    (C == 4'b1011) ? 7'b0000011 : // b
    (C == 4'b1100) ? 7'b1000110 : // c
    (C == 4'b1101) ? 7'b0100001 : // d
    (C == 4'b1110) ? 7'b0000110 : // e
    (C == 4'b1111) ? 7'b0001110 : // f
    7'b1111111; // blank

endmodule
